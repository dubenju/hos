conectix             �3�vpc   Wi2k    @      @  Z   ���\�,�6��h�jEL�                                                                                                                                                                                                                                                                                                                                                                                                                                            cxsparse��������             
    ���m                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ����������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        conectix             �3�vpc   Wi2k    @      @  Z   ���\�,�6��h�jEL�                                                                                                                                                                                                                                                                                                                                                                                                                                            